module TFF(T, Clock, Q);
input T, Clock;
output reg Q;

always@(posedge Clock)




