module count4bit(T, Clock, Q);
input T, Clock;
output reg Q;
//from textbook pg 298


endmodule
