 module lab8();
 