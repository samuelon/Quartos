//module lab8();
//endmodule