module FF(D,Clock,Q,Qn);
